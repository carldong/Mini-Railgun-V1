.SUBCKT OPA134   1 2 3 4 5
C1   11 12 3.240E-12
C2    6  7 8.000E-12
CSS  10 99 1.000E-30
DC    5 53 DX
DE   54  5 DX
DLP  90 91 DX
DLN  92 90 DX
DP    4  3 DX
EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
FB    7 99 POLY(5) VB VC VE VLP VLN 0 248.0E6 -250E6 250E6 250E6 -250E6
GA    6  0 11 12 402.0E-6
GCM   0  6 10 99 4.020E-9
ISS   3 10 DC 160.0E-6
HLIM 90  0 VLIM 1E3
J1   11  2 10 JX
J2   12  1 10 JX
R2    6  9 100.0E3
RD1   4 11 2.490E3
RD2   4 12 2.490E3
RO1   8  5 20
RO2   7 99 20
RP    3  4 7.500E3
RSS  10 99 1.250E6
VB    9  0 DC 0
VC    3 53 DC 1.200
VE   54  4 DC .9
VLIM  7  8 DC 0
VLP  91  0 DC 40
VLN   0 92 DC 40
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=2.500E-15 BETA=1.010E-3 VTO=-1)
.ENDS
V2 Vsig1 0 sin(0 5 500)
V1 3 0 DC 4.5V
R3 Vout1 0 1
R2 0 1 1K
R1 1 Vout1 10K
V3 2 0 DC -4.5V
XU1 Vsig1 1 3 2 Vout1 OPA134
.OP
.TRAN 50US 1.05S 1S
.PROBE V(Vsig1) V(Vout1)
.end
